��- -   C o d e   y o u r   t e s t b e n c h   h e r e  
 l i b r a r y   I E E E ;  
 u s e   I E E E . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 u s e   I E E E . n u m e r i c _ s t d . a l l ;  
  
 e n t i t y   k o l o _ t b   i s  
 	 g e n e r i c ( n   :   i n t e g e r   : =   4 ) ;  
 e n d   e n t i t y ;  
  
 a r c h i t e c t u r e   k o l o _ t b _ a r c h   o f   k o l o _ t b   i s  
 s i g n a l   A   ,   B   , D   :   s t d _ l o g i c _ v e c t o r ( n   d o w n t o   0 ) ;  
 s i g n a l   C   :   s t d _ l o g i c ;  
 b e g i n  
 	 D U T 1 : e n t i t y   w o r k . K o l o ( K o l o _ a r c h )  
         	 g e n e r i c   m a p ( n   = >   n )  
                 p o r t   m a p ( A   = >   A   ,   B = >   B   ,   D   = >   D   ,   C = >   C ) ;  
         S T I M U L U S :   p r o c e s s  
         	 b e g i n  
                 	 C   < =   ' 0 ' ;  
                 	 A   < =   " 1 0 1 0 0 " ;  
                         B   < =   " 0 0 0 0 0 " ;  
                         w a i t   f o r   2 0 0   n s ;  
         e n d   p r o c e s s ;  
 e n d   a r c h i t e c t u r e ;       