��- -   C o d e   y o u r   d e s i g n   h e r e  
 l i b r a r y   I E E E ;  
 u s e   I E E E . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 u s e   I E E E . n u m e r i c _ s t d . a l l ;  
  
 e n t i t y   O r G a t e   i s  
 	 p o r t ( A   :   i n   s t d _ l o g i c ;  
         	   B   :   i n   s t d _ l o g i c ;  
                   Y   :   o u t   s t d _ l o g i c ) ;  
 e n d   e n t i t y ;  
  
 a r c h i t e c t u r e   O r G a t e _ a r c h   o f   O r G a t e   i s  
 b e g i n  
 	 Y   < =   A   o r   B ;  
 e n d   a r c h i t e c t u r e ;  
  
 l i b r a r y   I E E E ;  
 u s e   I E E E . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 u s e   I E E E . n u m e r i c _ s t d . a l l ;  
  
 e n t i t y   X o r G a t e   i s  
 	 p o r t ( A   :   i n   s t d _ l o g i c ;  
         	   B   :   i n   s t d _ l o g i c ;  
                   Y   :   o u t   s t d _ l o g i c ) ;  
 e n d   e n t i t y ;  
  
 a r c h i t e c t u r e   X o r G a t e _ a r c h   o f   X o r G a t e   i s  
 b e g i n  
 	 Y   < =   A   x o r   B ;  
 e n d   a r c h i t e c t u r e ;  
  
  
  
 - -   S A D   I D E   O N O   P R A V O - -  
 l i b r a r y   I E E E ;  
 u s e   I E E E . s t d _ l o g i c _ 1 1 6 4 . a l l ;  
 u s e   I E E E . n u m e r i c _ s t d . a l l ;  
  
 e n t i t y   K o l o   i s  
 	 g e n e r i c ( n   :   i n t e g e r   : =   4 ) ;  
         p o r t ( A   :   i n   s t d _ l o g i c _ v e c t o r ( n   d o w n t o   0 ) ;  
         	   B   :   i n   s t d _ l o g i c _ v e c t o r ( n   d o w n t o   0 ) ;  
                   C   :   i n   s t d _ l o g i c ;  
                   D   :   o u t   s t d _ l o g i c _ v e c t o r ( n   d o w n t o   0 ) ) ;  
 e n d   e n t i t y ;  
  
 a r c h i t e c t u r e   K o l o _ a r c h   o f   K o l o   i s  
 s i g n a l   C _ u l a z   :   s t d _ l o g i c _ v e c t o r ( n   d o w n t o   0 ) ;  
 s i g n a l   X o r _ i z l a z   :   s t d _ l o g i c _ v e c t o r ( n   d o w n t o   0 ) ;  
 b e g i n  
 	 C _ u l a z ( 0 )   < =   C ;  
          
         F o r L b l   :   f o r   i   i n   0   t o   n   g e n e r a t e  
         b e g i n  
         	 I f 1 l b l   :   i f   i = 0   g e n e r a t e  
                 X o r _ G a t e :   e n t i t y   w o r k . X o r G a t e ( X o r G a t e _ a r c h )  
                 	 p o r t   m a p ( A   = >   A ( 0 )   ,   B   = >   B ( 0 )   ,   Y   = >   X o r _ i z l a z ( 0 ) ) ;  
                          
                 O r _ G a t e :   e n t i t y   w o r k . O r G a t e ( O r G a t e _ a r c h )  
                 	 p o r t   m a p ( A   = >   X o r _ i z l a z ( 0 )   ,   B   = >   C _ u l a z ( 0 )   ,   Y   = > D ( 0 ) ) ;  
                 C _ u l a z ( i + 1 )   < =   D ( 0 ) ;  
                 e n d   g e n e r a t e ;  
                  
                 I f 2 l b l   :   i f   i / = 0   a n d   i / = n   g e n e r a t e  
                 X o r _ G a t e   :   e n t i t y   w o r k . X o r G a t e ( X o r G a t e _ a r c h )  
                 	 p o r t   m a p ( A   = >   A ( i )   ,   B = >   B ( i )   ,   Y = > X o r _ i z l a z ( i ) ) ;  
                 O r _ G a t e :   e n t i t y   w o r k . O r G a t e ( O r G a t e _ a r c h )  
                 	 p o r t   m a p ( A   = >   X o r _ i z l a z ( i )   ,   B   = >   C _ u l a z ( i )   ,   Y   = > D ( i ) ) ;  
                 C _ u l a z ( i + 1 )   < =   D ( i ) ;  
                 e n d   g e n e r a t e ;  
                  
                   I f 3 l b l   :   i f   i = n   g e n e r a t e  
                 X o r _ G a t e   :   e n t i t y   w o r k . X o r G a t e ( X o r G a t e _ a r c h )  
                 	 p o r t   m a p ( A   = >   A ( i )   ,   B = >   B ( i )   ,   Y = > X o r _ i z l a z ( i ) ) ;  
                 O r _ G a t e :   e n t i t y   w o r k . O r G a t e ( O r G a t e _ a r c h )  
                 	 p o r t   m a p ( A   = >   X o r _ i z l a z ( i )   ,   B   = >   C _ u l a z ( i )   ,   Y   = > D ( i ) ) ;  
               e n d   g e n e r a t e ;  
                
         e n d   g e n e r a t e ;  
 e n d   a r c h i t e c t u r e ; 